`define DATA_WIDTH 16

