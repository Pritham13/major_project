module sync_fifo #(
    parameter DEPTH = 8,
    parameter type DTYPE = int
) (
    input        rstn,       // Active low reset
    input        clk,        // Clock
    input        fifo_wreq,  // Write enable
    input        fifo_rreq,  // Read enable
    input  DTYPE din,        // Data written into FIFO
    output DTYPE dout,       // Data read from FIFO
    output       empty,      // FIFO is empty when high
    output       full        // FIFO is full when high
);


  reg [$clog2(DEPTH)-1:0]   wptr;
  reg [$clog2(DEPTH)-1:0]   rptr;

  DTYPE    fifo[DEPTH];

  always @(posedge clk) begin
    if (!rstn) begin
      wptr <= 0;
    end else begin
      if (fifo_wreq & !full) begin
        fifo[wptr] <= din;
        wptr <= wptr + 1;
      end
    end
  end
  /*
  initial begin
    $monitor("[%0t] [FIFO] fifo_wreq=%0b din=0x%0h fifo_rreq=%0b dout=0x%0h empty=%0b full=%0b",
             $time, fifo_wreq, din, fifo_rreq, dout, empty, full);
  end
*/
  always @(posedge clk) begin
    if (!rstn) begin
      rptr <= 0;
    end else begin
      if (fifo_rreq & !empty) begin
        dout <= fifo[rptr];
        rptr <= rptr + 1;
      end
    end
  end

  assign full  = (wptr + 1) == rptr;
  assign empty = wptr == rptr;
endmodule
