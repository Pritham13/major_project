package fsm_pkg;
  
  // enums for request fsm 
  typedef enum {
    INITIAL_ST ,
    SAMPLE_DATA_ST,
    WRT_REQ_ST,
    WAIT_ST
    } req_states_e ;
endpackage
